// soc_system.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk_clk,                               //                       clk.clk
		input  wire        hps_0_f2h_cold_reset_req_reset_n,      //  hps_0_f2h_cold_reset_req.reset_n
		input  wire        hps_0_f2h_debug_reset_req_reset_n,     // hps_0_f2h_debug_reset_req.reset_n
		input  wire [27:0] hps_0_f2h_stm_hw_events_stm_hwevents,  //   hps_0_f2h_stm_hw_events.stm_hwevents
		input  wire        hps_0_f2h_warm_reset_req_reset_n,      //  hps_0_f2h_warm_reset_req.reset_n
		output wire        hps_0_h2f_reset_reset_n,               //           hps_0_h2f_reset.reset_n
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK, //              hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,   //                          .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,   //                          .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,   //                          .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,   //                          .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,   //                          .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,   //                          .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,    //                          .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL, //                          .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL, //                          .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK, //                          .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,   //                          .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,   //                          .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,   //                          .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,     //                          .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,      //                          .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,      //                          .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,     //                          .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,      //                          .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,      //                          .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,      //                          .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,      //                          .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,      //                          .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,      //                          .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,      //                          .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,      //                          .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,      //                          .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,      //                          .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,     //                          .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,     //                          .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,     //                          .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,     //                          .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,    //                          .hps_io_spim1_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,   //                          .hps_io_spim1_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,   //                          .hps_io_spim1_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,    //                          .hps_io_spim1_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,     //                          .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,     //                          .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,     //                          .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,     //                          .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,     //                          .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,     //                          .hps_io_i2c1_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,  //                          .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,  //                          .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,  //                          .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,  //                          .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,  //                          .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,  //                          .hps_io_gpio_inst_GPIO61
		inout  wire        i2c_avalon_bridge0_scl,                //        i2c_avalon_bridge0.scl
		inout  wire        i2c_avalon_bridge0_sda,                //                          .sda
		inout  wire        i2c_avalon_bridge1_scl,                //        i2c_avalon_bridge1.scl
		inout  wire        i2c_avalon_bridge1_sda,                //                          .sda
		output wire [14:0] memory_mem_a,                          //                    memory.mem_a
		output wire [2:0]  memory_mem_ba,                         //                          .mem_ba
		output wire        memory_mem_ck,                         //                          .mem_ck
		output wire        memory_mem_ck_n,                       //                          .mem_ck_n
		output wire        memory_mem_cke,                        //                          .mem_cke
		output wire        memory_mem_cs_n,                       //                          .mem_cs_n
		output wire        memory_mem_ras_n,                      //                          .mem_ras_n
		output wire        memory_mem_cas_n,                      //                          .mem_cas_n
		output wire        memory_mem_we_n,                       //                          .mem_we_n
		output wire        memory_mem_reset_n,                    //                          .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                         //                          .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                        //                          .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                      //                          .mem_dqs_n
		output wire        memory_mem_odt,                        //                          .mem_odt
		output wire [3:0]  memory_mem_dm,                         //                          .mem_dm
		input  wire        memory_oct_rzqin,                      //                          .oct_rzqin
		input  wire        reset_reset_n                          //                     reset.reset_n
	);

	wire    [1:0] hps_0_h2f_axi_master_awburst;                                     // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                       // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire    [7:0] hps_0_h2f_axi_master_wstrb;                                       // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_wready;                                      // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [11:0] hps_0_h2f_axi_master_rid;                                         // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_rready;                                      // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                       // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire   [11:0] hps_0_h2f_axi_master_wid;                                         // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                     // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire          hps_0_h2f_axi_master_wvalid;                                      // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                      // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                      // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                      // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire   [63:0] hps_0_h2f_axi_master_wdata;                                       // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_arvalid;                                     // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                     // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire   [11:0] hps_0_h2f_axi_master_arid;                                        // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                      // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                      // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                      // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                       // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire          hps_0_h2f_axi_master_arready;                                     // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire   [63:0] hps_0_h2f_axi_master_rdata;                                       // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire          hps_0_h2f_axi_master_awready;                                     // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                     // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                      // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire          hps_0_h2f_axi_master_bready;                                      // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire          hps_0_h2f_axi_master_rlast;                                       // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire          hps_0_h2f_axi_master_wlast;                                       // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                       // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire   [11:0] hps_0_h2f_axi_master_awid;                                        // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire   [11:0] hps_0_h2f_axi_master_bid;                                         // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire          hps_0_h2f_axi_master_bvalid;                                      // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                      // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire          hps_0_h2f_axi_master_awvalid;                                     // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire          hps_0_h2f_axi_master_rvalid;                                      // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire   [31:0] fpga_only_master_master_readdata;                                 // mm_interconnect_0:fpga_only_master_master_readdata -> fpga_only_master:master_readdata
	wire          fpga_only_master_master_waitrequest;                              // mm_interconnect_0:fpga_only_master_master_waitrequest -> fpga_only_master:master_waitrequest
	wire   [31:0] fpga_only_master_master_address;                                  // fpga_only_master:master_address -> mm_interconnect_0:fpga_only_master_master_address
	wire          fpga_only_master_master_read;                                     // fpga_only_master:master_read -> mm_interconnect_0:fpga_only_master_master_read
	wire    [3:0] fpga_only_master_master_byteenable;                               // fpga_only_master:master_byteenable -> mm_interconnect_0:fpga_only_master_master_byteenable
	wire          fpga_only_master_master_readdatavalid;                            // mm_interconnect_0:fpga_only_master_master_readdatavalid -> fpga_only_master:master_readdatavalid
	wire          fpga_only_master_master_write;                                    // fpga_only_master:master_write -> mm_interconnect_0:fpga_only_master_master_write
	wire   [31:0] fpga_only_master_master_writedata;                                // fpga_only_master:master_writedata -> mm_interconnect_0:fpga_only_master_master_writedata
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                                  // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                                    // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                                    // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_wready;                                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                                      // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_rready;                                   // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                                    // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                                      // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                                  // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire          hps_0_h2f_lw_axi_master_wvalid;                                   // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                                   // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                                   // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                                   // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                                    // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_arvalid;                                  // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                                  // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                                     // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                                   // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                                   // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                                   // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire          hps_0_h2f_lw_axi_master_arready;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire          hps_0_h2f_lw_axi_master_awready;                                  // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                                  // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                                   // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire          hps_0_h2f_lw_axi_master_bready;                                   // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire          hps_0_h2f_lw_axi_master_rlast;                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire          hps_0_h2f_lw_axi_master_wlast;                                    // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                                    // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                                     // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                                      // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire          hps_0_h2f_lw_axi_master_bvalid;                                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                                   // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire          hps_0_h2f_lw_axi_master_awvalid;                                  // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire          hps_0_h2f_lw_axi_master_rvalid;                                   // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire          mm_interconnect_0_onchip_memory2_0_s1_chipselect;                 // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire   [63:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                   // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [12:0] mm_interconnect_0_onchip_memory2_0_s1_address;                    // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire    [7:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                 // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire          mm_interconnect_0_onchip_memory2_0_s1_write;                      // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire   [63:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                  // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire          mm_interconnect_0_onchip_memory2_0_s1_clken;                      // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;           // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;        // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;              // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [31:0] mm_interconnect_0_intr_capturer_0_avalon_slave_0_readdata;        // intr_capturer_0:rddata -> mm_interconnect_0:intr_capturer_0_avalon_slave_0_readdata
	wire    [0:0] mm_interconnect_0_intr_capturer_0_avalon_slave_0_address;         // mm_interconnect_0:intr_capturer_0_avalon_slave_0_address -> intr_capturer_0:addr
	wire          mm_interconnect_0_intr_capturer_0_avalon_slave_0_read;            // mm_interconnect_0:intr_capturer_0_avalon_slave_0_read -> intr_capturer_0:read
	wire   [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;              // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire    [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;               // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire   [31:0] mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_readdata;    // I2C_avalon_bridge_0:readdata -> mm_interconnect_0:I2C_avalon_bridge_0_avalon_slave_0_readdata
	wire          mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_waitrequest; // I2C_avalon_bridge_0:waitrequest -> mm_interconnect_0:I2C_avalon_bridge_0_avalon_slave_0_waitrequest
	wire    [2:0] mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_address;     // mm_interconnect_0:I2C_avalon_bridge_0_avalon_slave_0_address -> I2C_avalon_bridge_0:address
	wire          mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_read;        // mm_interconnect_0:I2C_avalon_bridge_0_avalon_slave_0_read -> I2C_avalon_bridge_0:read
	wire          mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_write;       // mm_interconnect_0:I2C_avalon_bridge_0_avalon_slave_0_write -> I2C_avalon_bridge_0:write
	wire   [31:0] mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_writedata;   // mm_interconnect_0:I2C_avalon_bridge_0_avalon_slave_0_writedata -> I2C_avalon_bridge_0:writedata
	wire   [31:0] mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_readdata;    // I2C_avalon_bridge_1:readdata -> mm_interconnect_0:I2C_avalon_bridge_1_avalon_slave_0_readdata
	wire          mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_waitrequest; // I2C_avalon_bridge_1:waitrequest -> mm_interconnect_0:I2C_avalon_bridge_1_avalon_slave_0_waitrequest
	wire    [2:0] mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_address;     // mm_interconnect_0:I2C_avalon_bridge_1_avalon_slave_0_address -> I2C_avalon_bridge_1:address
	wire          mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_read;        // mm_interconnect_0:I2C_avalon_bridge_1_avalon_slave_0_read -> I2C_avalon_bridge_1:read
	wire          mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_write;       // mm_interconnect_0:I2C_avalon_bridge_1_avalon_slave_0_write -> I2C_avalon_bridge_1:write
	wire   [31:0] mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_writedata;   // mm_interconnect_0:I2C_avalon_bridge_1_avalon_slave_0_writedata -> I2C_avalon_bridge_1:writedata
	wire   [31:0] hps_only_master_master_readdata;                                  // mm_interconnect_1:hps_only_master_master_readdata -> hps_only_master:master_readdata
	wire          hps_only_master_master_waitrequest;                               // mm_interconnect_1:hps_only_master_master_waitrequest -> hps_only_master:master_waitrequest
	wire   [31:0] hps_only_master_master_address;                                   // hps_only_master:master_address -> mm_interconnect_1:hps_only_master_master_address
	wire          hps_only_master_master_read;                                      // hps_only_master:master_read -> mm_interconnect_1:hps_only_master_master_read
	wire    [3:0] hps_only_master_master_byteenable;                                // hps_only_master:master_byteenable -> mm_interconnect_1:hps_only_master_master_byteenable
	wire          hps_only_master_master_readdatavalid;                             // mm_interconnect_1:hps_only_master_master_readdatavalid -> hps_only_master:master_readdatavalid
	wire          hps_only_master_master_write;                                     // hps_only_master:master_write -> mm_interconnect_1:hps_only_master_master_write
	wire   [31:0] hps_only_master_master_writedata;                                 // hps_only_master:master_writedata -> mm_interconnect_1:hps_only_master_master_writedata
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_awburst;                    // mm_interconnect_1:hps_0_f2h_axi_slave_awburst -> hps_0:f2h_AWBURST
	wire    [4:0] mm_interconnect_1_hps_0_f2h_axi_slave_awuser;                     // mm_interconnect_1:hps_0_f2h_axi_slave_awuser -> hps_0:f2h_AWUSER
	wire    [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_arlen;                      // mm_interconnect_1:hps_0_f2h_axi_slave_arlen -> hps_0:f2h_ARLEN
	wire   [15:0] mm_interconnect_1_hps_0_f2h_axi_slave_wstrb;                      // mm_interconnect_1:hps_0_f2h_axi_slave_wstrb -> hps_0:f2h_WSTRB
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_wready;                     // hps_0:f2h_WREADY -> mm_interconnect_1:hps_0_f2h_axi_slave_wready
	wire    [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_rid;                        // hps_0:f2h_RID -> mm_interconnect_1:hps_0_f2h_axi_slave_rid
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_rready;                     // mm_interconnect_1:hps_0_f2h_axi_slave_rready -> hps_0:f2h_RREADY
	wire    [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_awlen;                      // mm_interconnect_1:hps_0_f2h_axi_slave_awlen -> hps_0:f2h_AWLEN
	wire    [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_wid;                        // mm_interconnect_1:hps_0_f2h_axi_slave_wid -> hps_0:f2h_WID
	wire    [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_arcache;                    // mm_interconnect_1:hps_0_f2h_axi_slave_arcache -> hps_0:f2h_ARCACHE
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_wvalid;                     // mm_interconnect_1:hps_0_f2h_axi_slave_wvalid -> hps_0:f2h_WVALID
	wire   [31:0] mm_interconnect_1_hps_0_f2h_axi_slave_araddr;                     // mm_interconnect_1:hps_0_f2h_axi_slave_araddr -> hps_0:f2h_ARADDR
	wire    [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_arprot;                     // mm_interconnect_1:hps_0_f2h_axi_slave_arprot -> hps_0:f2h_ARPROT
	wire    [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_awprot;                     // mm_interconnect_1:hps_0_f2h_axi_slave_awprot -> hps_0:f2h_AWPROT
	wire  [127:0] mm_interconnect_1_hps_0_f2h_axi_slave_wdata;                      // mm_interconnect_1:hps_0_f2h_axi_slave_wdata -> hps_0:f2h_WDATA
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_arvalid;                    // mm_interconnect_1:hps_0_f2h_axi_slave_arvalid -> hps_0:f2h_ARVALID
	wire    [3:0] mm_interconnect_1_hps_0_f2h_axi_slave_awcache;                    // mm_interconnect_1:hps_0_f2h_axi_slave_awcache -> hps_0:f2h_AWCACHE
	wire    [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_arid;                       // mm_interconnect_1:hps_0_f2h_axi_slave_arid -> hps_0:f2h_ARID
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_arlock;                     // mm_interconnect_1:hps_0_f2h_axi_slave_arlock -> hps_0:f2h_ARLOCK
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_awlock;                     // mm_interconnect_1:hps_0_f2h_axi_slave_awlock -> hps_0:f2h_AWLOCK
	wire   [31:0] mm_interconnect_1_hps_0_f2h_axi_slave_awaddr;                     // mm_interconnect_1:hps_0_f2h_axi_slave_awaddr -> hps_0:f2h_AWADDR
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_bresp;                      // hps_0:f2h_BRESP -> mm_interconnect_1:hps_0_f2h_axi_slave_bresp
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_arready;                    // hps_0:f2h_ARREADY -> mm_interconnect_1:hps_0_f2h_axi_slave_arready
	wire  [127:0] mm_interconnect_1_hps_0_f2h_axi_slave_rdata;                      // hps_0:f2h_RDATA -> mm_interconnect_1:hps_0_f2h_axi_slave_rdata
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_awready;                    // hps_0:f2h_AWREADY -> mm_interconnect_1:hps_0_f2h_axi_slave_awready
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_arburst;                    // mm_interconnect_1:hps_0_f2h_axi_slave_arburst -> hps_0:f2h_ARBURST
	wire    [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_arsize;                     // mm_interconnect_1:hps_0_f2h_axi_slave_arsize -> hps_0:f2h_ARSIZE
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_bready;                     // mm_interconnect_1:hps_0_f2h_axi_slave_bready -> hps_0:f2h_BREADY
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_rlast;                      // hps_0:f2h_RLAST -> mm_interconnect_1:hps_0_f2h_axi_slave_rlast
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_wlast;                      // mm_interconnect_1:hps_0_f2h_axi_slave_wlast -> hps_0:f2h_WLAST
	wire    [1:0] mm_interconnect_1_hps_0_f2h_axi_slave_rresp;                      // hps_0:f2h_RRESP -> mm_interconnect_1:hps_0_f2h_axi_slave_rresp
	wire    [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_awid;                       // mm_interconnect_1:hps_0_f2h_axi_slave_awid -> hps_0:f2h_AWID
	wire    [7:0] mm_interconnect_1_hps_0_f2h_axi_slave_bid;                        // hps_0:f2h_BID -> mm_interconnect_1:hps_0_f2h_axi_slave_bid
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_bvalid;                     // hps_0:f2h_BVALID -> mm_interconnect_1:hps_0_f2h_axi_slave_bvalid
	wire    [2:0] mm_interconnect_1_hps_0_f2h_axi_slave_awsize;                     // mm_interconnect_1:hps_0_f2h_axi_slave_awsize -> hps_0:f2h_AWSIZE
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_awvalid;                    // mm_interconnect_1:hps_0_f2h_axi_slave_awvalid -> hps_0:f2h_AWVALID
	wire    [4:0] mm_interconnect_1_hps_0_f2h_axi_slave_aruser;                     // mm_interconnect_1:hps_0_f2h_axi_slave_aruser -> hps_0:f2h_ARUSER
	wire          mm_interconnect_1_hps_0_f2h_axi_slave_rvalid;                     // hps_0:f2h_RVALID -> mm_interconnect_1:hps_0_f2h_axi_slave_rvalid
	wire   [31:0] hps_0_f2h_irq0_irq;                                               // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                               // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire   [31:0] intr_capturer_0_interrupt_receiver_irq;                           // irq_mapper_002:sender_irq -> intr_capturer_0:interrupt_in
	wire          irq_mapper_receiver0_irq;                                         // jtag_uart:av_irq -> [irq_mapper:receiver0_irq, irq_mapper_002:receiver0_irq]
	wire          rst_controller_reset_out_reset;                                   // rst_controller:reset_out -> [I2C_avalon_bridge_0:reset, I2C_avalon_bridge_1:reset, intr_capturer_0:rst_n, irq_mapper_002:reset, jtag_uart:rst_n, mm_interconnect_0:fpga_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:onchip_memory2_0_reset1_reset_bridge_in_reset_reset, mm_interconnect_1:hps_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_only_master_master_translator_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_translator:in_reset, sysid_qsys:reset_n]
	wire          rst_controller_reset_out_reset_req;                               // rst_controller:reset_req -> [onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                               // rst_controller_001:reset_out -> [mm_interconnect_0:hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset]

	I2C_avalon_bridge i2c_avalon_bridge_0 (
		.reset       (rst_controller_reset_out_reset),                                   //          reset.reset
		.address     (mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_address),     // avalon_slave_0.address
		.write       (mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_write),       //               .write
		.writedata   (mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_writedata),   //               .writedata
		.read        (mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_read),        //               .read
		.readdata    (mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_readdata),    //               .readdata
		.waitrequest (mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_waitrequest), //               .waitrequest
		.scl         (i2c_avalon_bridge0_scl),                                           //    conduit_end.scl
		.sda         (i2c_avalon_bridge0_sda),                                           //               .sda
		.clock       (clk_clk)                                                           //     clock_sink.clk
	);

	I2C_avalon_bridge i2c_avalon_bridge_1 (
		.reset       (rst_controller_reset_out_reset),                                   //          reset.reset
		.address     (mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_address),     // avalon_slave_0.address
		.write       (mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_write),       //               .write
		.writedata   (mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_writedata),   //               .writedata
		.read        (mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_read),        //               .read
		.readdata    (mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_readdata),    //               .readdata
		.waitrequest (mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_waitrequest), //               .waitrequest
		.scl         (i2c_avalon_bridge1_scl),                                           //    conduit_end.scl
		.sda         (i2c_avalon_bridge1_sda),                                           //               .sda
		.clock       (clk_clk)                                                           //     clock_sink.clk
	);

	soc_system_fpga_only_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) fpga_only_master (
		.clk_clk              (clk_clk),                               //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                        //    clk_reset.reset
		.master_address       (fpga_only_master_master_address),       //       master.address
		.master_readdata      (fpga_only_master_master_readdata),      //             .readdata
		.master_read          (fpga_only_master_master_read),          //             .read
		.master_write         (fpga_only_master_master_write),         //             .write
		.master_writedata     (fpga_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (fpga_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (fpga_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (fpga_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                       // master_reset.reset
	);

	soc_system_hps_0 #(
		.F2S_Width (3),
		.S2F_Width (2)
	) hps_0 (
		.f2h_cold_rst_req_n       (hps_0_f2h_cold_reset_req_reset_n),              //  f2h_cold_reset_req.reset_n
		.f2h_dbg_rst_req_n        (hps_0_f2h_debug_reset_req_reset_n),             // f2h_debug_reset_req.reset_n
		.f2h_warm_rst_req_n       (hps_0_f2h_warm_reset_req_reset_n),              //  f2h_warm_reset_req.reset_n
		.f2h_stm_hwevents         (hps_0_f2h_stm_hw_events_stm_hwevents),          //   f2h_stm_hw_events.stm_hwevents
		.mem_a                    (memory_mem_a),                                  //              memory.mem_a
		.mem_ba                   (memory_mem_ba),                                 //                    .mem_ba
		.mem_ck                   (memory_mem_ck),                                 //                    .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                               //                    .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                //                    .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                               //                    .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                              //                    .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                              //                    .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                               //                    .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                            //                    .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                 //                    .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                //                    .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                              //                    .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                //                    .mem_odt
		.mem_dm                   (memory_mem_dm),                                 //                    .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                              //                    .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_hps_io_hps_io_emac1_inst_TX_CLK),         //              hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_hps_io_hps_io_emac1_inst_TXD0),           //                    .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_hps_io_hps_io_emac1_inst_TXD1),           //                    .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_hps_io_hps_io_emac1_inst_TXD2),           //                    .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_hps_io_hps_io_emac1_inst_TXD3),           //                    .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_hps_io_hps_io_emac1_inst_RXD0),           //                    .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_hps_io_hps_io_emac1_inst_MDIO),           //                    .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_hps_io_hps_io_emac1_inst_MDC),            //                    .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_hps_io_hps_io_emac1_inst_RX_CTL),         //                    .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_hps_io_hps_io_emac1_inst_TX_CTL),         //                    .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_hps_io_hps_io_emac1_inst_RX_CLK),         //                    .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_hps_io_hps_io_emac1_inst_RXD1),           //                    .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_hps_io_hps_io_emac1_inst_RXD2),           //                    .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_hps_io_hps_io_emac1_inst_RXD3),           //                    .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_0_hps_io_hps_io_sdio_inst_CMD),             //                    .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_hps_io_hps_io_sdio_inst_D0),              //                    .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_hps_io_hps_io_sdio_inst_D1),              //                    .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_hps_io_hps_io_sdio_inst_CLK),             //                    .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_hps_io_hps_io_sdio_inst_D2),              //                    .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_hps_io_hps_io_sdio_inst_D3),              //                    .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_hps_io_hps_io_usb1_inst_D0),              //                    .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_hps_io_hps_io_usb1_inst_D1),              //                    .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_hps_io_hps_io_usb1_inst_D2),              //                    .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_hps_io_hps_io_usb1_inst_D3),              //                    .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_hps_io_hps_io_usb1_inst_D4),              //                    .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_hps_io_hps_io_usb1_inst_D5),              //                    .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_hps_io_hps_io_usb1_inst_D6),              //                    .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_hps_io_hps_io_usb1_inst_D7),              //                    .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_hps_io_hps_io_usb1_inst_CLK),             //                    .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_hps_io_hps_io_usb1_inst_STP),             //                    .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_hps_io_hps_io_usb1_inst_DIR),             //                    .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_hps_io_hps_io_usb1_inst_NXT),             //                    .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_0_hps_io_hps_io_spim1_inst_CLK),            //                    .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_0_hps_io_hps_io_spim1_inst_MOSI),           //                    .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_0_hps_io_hps_io_spim1_inst_MISO),           //                    .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_0_hps_io_hps_io_spim1_inst_SS0),            //                    .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_0_hps_io_hps_io_uart0_inst_RX),             //                    .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_hps_io_hps_io_uart0_inst_TX),             //                    .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_hps_io_hps_io_i2c0_inst_SDA),             //                    .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_hps_io_hps_io_i2c0_inst_SCL),             //                    .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_0_hps_io_hps_io_i2c1_inst_SDA),             //                    .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_0_hps_io_hps_io_i2c1_inst_SCL),             //                    .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_0_hps_io_hps_io_gpio_inst_GPIO09),          //                    .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_0_hps_io_hps_io_gpio_inst_GPIO35),          //                    .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_0_hps_io_hps_io_gpio_inst_GPIO40),          //                    .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO53  (hps_0_hps_io_hps_io_gpio_inst_GPIO53),          //                    .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_0_hps_io_hps_io_gpio_inst_GPIO54),          //                    .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_0_hps_io_hps_io_gpio_inst_GPIO61),          //                    .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),                       //           h2f_reset.reset_n
		.h2f_axi_clk              (clk_clk),                                       //       h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),                     //      h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),                   //                    .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),                    //                    .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),                   //                    .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),                  //                    .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),                   //                    .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),                  //                    .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),                   //                    .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),                  //                    .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),                  //                    .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),                      //                    .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),                    //                    .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),                    //                    .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),                    //                    .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),                   //                    .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),                   //                    .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),                      //                    .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),                    //                    .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),                   //                    .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),                   //                    .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),                     //                    .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),                   //                    .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),                    //                    .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),                   //                    .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),                  //                    .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),                   //                    .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),                  //                    .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),                   //                    .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),                  //                    .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),                  //                    .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),                      //                    .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),                    //                    .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),                    //                    .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),                    //                    .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),                   //                    .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),                   //                    .rready
		.f2h_axi_clk              (clk_clk),                                       //       f2h_axi_clock.clk
		.f2h_AWID                 (mm_interconnect_1_hps_0_f2h_axi_slave_awid),    //       f2h_axi_slave.awid
		.f2h_AWADDR               (mm_interconnect_1_hps_0_f2h_axi_slave_awaddr),  //                    .awaddr
		.f2h_AWLEN                (mm_interconnect_1_hps_0_f2h_axi_slave_awlen),   //                    .awlen
		.f2h_AWSIZE               (mm_interconnect_1_hps_0_f2h_axi_slave_awsize),  //                    .awsize
		.f2h_AWBURST              (mm_interconnect_1_hps_0_f2h_axi_slave_awburst), //                    .awburst
		.f2h_AWLOCK               (mm_interconnect_1_hps_0_f2h_axi_slave_awlock),  //                    .awlock
		.f2h_AWCACHE              (mm_interconnect_1_hps_0_f2h_axi_slave_awcache), //                    .awcache
		.f2h_AWPROT               (mm_interconnect_1_hps_0_f2h_axi_slave_awprot),  //                    .awprot
		.f2h_AWVALID              (mm_interconnect_1_hps_0_f2h_axi_slave_awvalid), //                    .awvalid
		.f2h_AWREADY              (mm_interconnect_1_hps_0_f2h_axi_slave_awready), //                    .awready
		.f2h_AWUSER               (mm_interconnect_1_hps_0_f2h_axi_slave_awuser),  //                    .awuser
		.f2h_WID                  (mm_interconnect_1_hps_0_f2h_axi_slave_wid),     //                    .wid
		.f2h_WDATA                (mm_interconnect_1_hps_0_f2h_axi_slave_wdata),   //                    .wdata
		.f2h_WSTRB                (mm_interconnect_1_hps_0_f2h_axi_slave_wstrb),   //                    .wstrb
		.f2h_WLAST                (mm_interconnect_1_hps_0_f2h_axi_slave_wlast),   //                    .wlast
		.f2h_WVALID               (mm_interconnect_1_hps_0_f2h_axi_slave_wvalid),  //                    .wvalid
		.f2h_WREADY               (mm_interconnect_1_hps_0_f2h_axi_slave_wready),  //                    .wready
		.f2h_BID                  (mm_interconnect_1_hps_0_f2h_axi_slave_bid),     //                    .bid
		.f2h_BRESP                (mm_interconnect_1_hps_0_f2h_axi_slave_bresp),   //                    .bresp
		.f2h_BVALID               (mm_interconnect_1_hps_0_f2h_axi_slave_bvalid),  //                    .bvalid
		.f2h_BREADY               (mm_interconnect_1_hps_0_f2h_axi_slave_bready),  //                    .bready
		.f2h_ARID                 (mm_interconnect_1_hps_0_f2h_axi_slave_arid),    //                    .arid
		.f2h_ARADDR               (mm_interconnect_1_hps_0_f2h_axi_slave_araddr),  //                    .araddr
		.f2h_ARLEN                (mm_interconnect_1_hps_0_f2h_axi_slave_arlen),   //                    .arlen
		.f2h_ARSIZE               (mm_interconnect_1_hps_0_f2h_axi_slave_arsize),  //                    .arsize
		.f2h_ARBURST              (mm_interconnect_1_hps_0_f2h_axi_slave_arburst), //                    .arburst
		.f2h_ARLOCK               (mm_interconnect_1_hps_0_f2h_axi_slave_arlock),  //                    .arlock
		.f2h_ARCACHE              (mm_interconnect_1_hps_0_f2h_axi_slave_arcache), //                    .arcache
		.f2h_ARPROT               (mm_interconnect_1_hps_0_f2h_axi_slave_arprot),  //                    .arprot
		.f2h_ARVALID              (mm_interconnect_1_hps_0_f2h_axi_slave_arvalid), //                    .arvalid
		.f2h_ARREADY              (mm_interconnect_1_hps_0_f2h_axi_slave_arready), //                    .arready
		.f2h_ARUSER               (mm_interconnect_1_hps_0_f2h_axi_slave_aruser),  //                    .aruser
		.f2h_RID                  (mm_interconnect_1_hps_0_f2h_axi_slave_rid),     //                    .rid
		.f2h_RDATA                (mm_interconnect_1_hps_0_f2h_axi_slave_rdata),   //                    .rdata
		.f2h_RRESP                (mm_interconnect_1_hps_0_f2h_axi_slave_rresp),   //                    .rresp
		.f2h_RLAST                (mm_interconnect_1_hps_0_f2h_axi_slave_rlast),   //                    .rlast
		.f2h_RVALID               (mm_interconnect_1_hps_0_f2h_axi_slave_rvalid),  //                    .rvalid
		.f2h_RREADY               (mm_interconnect_1_hps_0_f2h_axi_slave_rready),  //                    .rready
		.h2f_lw_axi_clk           (clk_clk),                                       //    h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                  //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                //                    .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                 //                    .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                //                    .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),               //                    .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                //                    .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),               //                    .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                //                    .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),               //                    .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),               //                    .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                   //                    .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                 //                    .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                 //                    .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                 //                    .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                //                    .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                //                    .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                   //                    .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                 //                    .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                //                    .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                //                    .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                  //                    .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                //                    .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                 //                    .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                //                    .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),               //                    .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                //                    .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),               //                    .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                //                    .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),               //                    .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),               //                    .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                   //                    .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                 //                    .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                 //                    .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                 //                    .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                //                    .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),                //                    .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                            //            f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                             //            f2h_irq1.irq
	);

	soc_system_fpga_only_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) hps_only_master (
		.clk_clk              (clk_clk),                              //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                       //    clk_reset.reset
		.master_address       (hps_only_master_master_address),       //       master.address
		.master_readdata      (hps_only_master_master_readdata),      //             .readdata
		.master_read          (hps_only_master_master_read),          //             .read
		.master_write         (hps_only_master_master_write),         //             .write
		.master_writedata     (hps_only_master_master_writedata),     //             .writedata
		.master_waitrequest   (hps_only_master_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (hps_only_master_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (hps_only_master_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                      // master_reset.reset
	);

	intr_capturer #(
		.NUM_INTR (32)
	) intr_capturer_0 (
		.clk          (clk_clk),                                                   //              clock.clk
		.rst_n        (~rst_controller_reset_out_reset),                           //         reset_sink.reset_n
		.addr         (mm_interconnect_0_intr_capturer_0_avalon_slave_0_address),  //     avalon_slave_0.address
		.read         (mm_interconnect_0_intr_capturer_0_avalon_slave_0_read),     //                   .read
		.rddata       (mm_interconnect_0_intr_capturer_0_avalon_slave_0_readdata), //                   .readdata
		.interrupt_in (intr_capturer_0_interrupt_receiver_irq)                     // interrupt_receiver.irq
	);

	soc_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	soc_system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	soc_system_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                        (hps_0_h2f_axi_master_awid),                                        //                                       hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                      (hps_0_h2f_axi_master_awaddr),                                      //                                                           .awaddr
		.hps_0_h2f_axi_master_awlen                                       (hps_0_h2f_axi_master_awlen),                                       //                                                           .awlen
		.hps_0_h2f_axi_master_awsize                                      (hps_0_h2f_axi_master_awsize),                                      //                                                           .awsize
		.hps_0_h2f_axi_master_awburst                                     (hps_0_h2f_axi_master_awburst),                                     //                                                           .awburst
		.hps_0_h2f_axi_master_awlock                                      (hps_0_h2f_axi_master_awlock),                                      //                                                           .awlock
		.hps_0_h2f_axi_master_awcache                                     (hps_0_h2f_axi_master_awcache),                                     //                                                           .awcache
		.hps_0_h2f_axi_master_awprot                                      (hps_0_h2f_axi_master_awprot),                                      //                                                           .awprot
		.hps_0_h2f_axi_master_awvalid                                     (hps_0_h2f_axi_master_awvalid),                                     //                                                           .awvalid
		.hps_0_h2f_axi_master_awready                                     (hps_0_h2f_axi_master_awready),                                     //                                                           .awready
		.hps_0_h2f_axi_master_wid                                         (hps_0_h2f_axi_master_wid),                                         //                                                           .wid
		.hps_0_h2f_axi_master_wdata                                       (hps_0_h2f_axi_master_wdata),                                       //                                                           .wdata
		.hps_0_h2f_axi_master_wstrb                                       (hps_0_h2f_axi_master_wstrb),                                       //                                                           .wstrb
		.hps_0_h2f_axi_master_wlast                                       (hps_0_h2f_axi_master_wlast),                                       //                                                           .wlast
		.hps_0_h2f_axi_master_wvalid                                      (hps_0_h2f_axi_master_wvalid),                                      //                                                           .wvalid
		.hps_0_h2f_axi_master_wready                                      (hps_0_h2f_axi_master_wready),                                      //                                                           .wready
		.hps_0_h2f_axi_master_bid                                         (hps_0_h2f_axi_master_bid),                                         //                                                           .bid
		.hps_0_h2f_axi_master_bresp                                       (hps_0_h2f_axi_master_bresp),                                       //                                                           .bresp
		.hps_0_h2f_axi_master_bvalid                                      (hps_0_h2f_axi_master_bvalid),                                      //                                                           .bvalid
		.hps_0_h2f_axi_master_bready                                      (hps_0_h2f_axi_master_bready),                                      //                                                           .bready
		.hps_0_h2f_axi_master_arid                                        (hps_0_h2f_axi_master_arid),                                        //                                                           .arid
		.hps_0_h2f_axi_master_araddr                                      (hps_0_h2f_axi_master_araddr),                                      //                                                           .araddr
		.hps_0_h2f_axi_master_arlen                                       (hps_0_h2f_axi_master_arlen),                                       //                                                           .arlen
		.hps_0_h2f_axi_master_arsize                                      (hps_0_h2f_axi_master_arsize),                                      //                                                           .arsize
		.hps_0_h2f_axi_master_arburst                                     (hps_0_h2f_axi_master_arburst),                                     //                                                           .arburst
		.hps_0_h2f_axi_master_arlock                                      (hps_0_h2f_axi_master_arlock),                                      //                                                           .arlock
		.hps_0_h2f_axi_master_arcache                                     (hps_0_h2f_axi_master_arcache),                                     //                                                           .arcache
		.hps_0_h2f_axi_master_arprot                                      (hps_0_h2f_axi_master_arprot),                                      //                                                           .arprot
		.hps_0_h2f_axi_master_arvalid                                     (hps_0_h2f_axi_master_arvalid),                                     //                                                           .arvalid
		.hps_0_h2f_axi_master_arready                                     (hps_0_h2f_axi_master_arready),                                     //                                                           .arready
		.hps_0_h2f_axi_master_rid                                         (hps_0_h2f_axi_master_rid),                                         //                                                           .rid
		.hps_0_h2f_axi_master_rdata                                       (hps_0_h2f_axi_master_rdata),                                       //                                                           .rdata
		.hps_0_h2f_axi_master_rresp                                       (hps_0_h2f_axi_master_rresp),                                       //                                                           .rresp
		.hps_0_h2f_axi_master_rlast                                       (hps_0_h2f_axi_master_rlast),                                       //                                                           .rlast
		.hps_0_h2f_axi_master_rvalid                                      (hps_0_h2f_axi_master_rvalid),                                      //                                                           .rvalid
		.hps_0_h2f_axi_master_rready                                      (hps_0_h2f_axi_master_rready),                                      //                                                           .rready
		.hps_0_h2f_lw_axi_master_awid                                     (hps_0_h2f_lw_axi_master_awid),                                     //                                    hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                   (hps_0_h2f_lw_axi_master_awaddr),                                   //                                                           .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                    (hps_0_h2f_lw_axi_master_awlen),                                    //                                                           .awlen
		.hps_0_h2f_lw_axi_master_awsize                                   (hps_0_h2f_lw_axi_master_awsize),                                   //                                                           .awsize
		.hps_0_h2f_lw_axi_master_awburst                                  (hps_0_h2f_lw_axi_master_awburst),                                  //                                                           .awburst
		.hps_0_h2f_lw_axi_master_awlock                                   (hps_0_h2f_lw_axi_master_awlock),                                   //                                                           .awlock
		.hps_0_h2f_lw_axi_master_awcache                                  (hps_0_h2f_lw_axi_master_awcache),                                  //                                                           .awcache
		.hps_0_h2f_lw_axi_master_awprot                                   (hps_0_h2f_lw_axi_master_awprot),                                   //                                                           .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                  (hps_0_h2f_lw_axi_master_awvalid),                                  //                                                           .awvalid
		.hps_0_h2f_lw_axi_master_awready                                  (hps_0_h2f_lw_axi_master_awready),                                  //                                                           .awready
		.hps_0_h2f_lw_axi_master_wid                                      (hps_0_h2f_lw_axi_master_wid),                                      //                                                           .wid
		.hps_0_h2f_lw_axi_master_wdata                                    (hps_0_h2f_lw_axi_master_wdata),                                    //                                                           .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                    (hps_0_h2f_lw_axi_master_wstrb),                                    //                                                           .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                    (hps_0_h2f_lw_axi_master_wlast),                                    //                                                           .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                   (hps_0_h2f_lw_axi_master_wvalid),                                   //                                                           .wvalid
		.hps_0_h2f_lw_axi_master_wready                                   (hps_0_h2f_lw_axi_master_wready),                                   //                                                           .wready
		.hps_0_h2f_lw_axi_master_bid                                      (hps_0_h2f_lw_axi_master_bid),                                      //                                                           .bid
		.hps_0_h2f_lw_axi_master_bresp                                    (hps_0_h2f_lw_axi_master_bresp),                                    //                                                           .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                   (hps_0_h2f_lw_axi_master_bvalid),                                   //                                                           .bvalid
		.hps_0_h2f_lw_axi_master_bready                                   (hps_0_h2f_lw_axi_master_bready),                                   //                                                           .bready
		.hps_0_h2f_lw_axi_master_arid                                     (hps_0_h2f_lw_axi_master_arid),                                     //                                                           .arid
		.hps_0_h2f_lw_axi_master_araddr                                   (hps_0_h2f_lw_axi_master_araddr),                                   //                                                           .araddr
		.hps_0_h2f_lw_axi_master_arlen                                    (hps_0_h2f_lw_axi_master_arlen),                                    //                                                           .arlen
		.hps_0_h2f_lw_axi_master_arsize                                   (hps_0_h2f_lw_axi_master_arsize),                                   //                                                           .arsize
		.hps_0_h2f_lw_axi_master_arburst                                  (hps_0_h2f_lw_axi_master_arburst),                                  //                                                           .arburst
		.hps_0_h2f_lw_axi_master_arlock                                   (hps_0_h2f_lw_axi_master_arlock),                                   //                                                           .arlock
		.hps_0_h2f_lw_axi_master_arcache                                  (hps_0_h2f_lw_axi_master_arcache),                                  //                                                           .arcache
		.hps_0_h2f_lw_axi_master_arprot                                   (hps_0_h2f_lw_axi_master_arprot),                                   //                                                           .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                  (hps_0_h2f_lw_axi_master_arvalid),                                  //                                                           .arvalid
		.hps_0_h2f_lw_axi_master_arready                                  (hps_0_h2f_lw_axi_master_arready),                                  //                                                           .arready
		.hps_0_h2f_lw_axi_master_rid                                      (hps_0_h2f_lw_axi_master_rid),                                      //                                                           .rid
		.hps_0_h2f_lw_axi_master_rdata                                    (hps_0_h2f_lw_axi_master_rdata),                                    //                                                           .rdata
		.hps_0_h2f_lw_axi_master_rresp                                    (hps_0_h2f_lw_axi_master_rresp),                                    //                                                           .rresp
		.hps_0_h2f_lw_axi_master_rlast                                    (hps_0_h2f_lw_axi_master_rlast),                                    //                                                           .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                   (hps_0_h2f_lw_axi_master_rvalid),                                   //                                                           .rvalid
		.hps_0_h2f_lw_axi_master_rready                                   (hps_0_h2f_lw_axi_master_rready),                                   //                                                           .rready
		.clk_0_clk_clk                                                    (clk_clk),                                                          //                                                  clk_0_clk.clk
		.fpga_only_master_clk_reset_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                                   //           fpga_only_master_clk_reset_reset_bridge_in_reset.reset
		.hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                               // hps_0_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.onchip_memory2_0_reset1_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),                                   //              onchip_memory2_0_reset1_reset_bridge_in_reset.reset
		.fpga_only_master_master_address                                  (fpga_only_master_master_address),                                  //                                    fpga_only_master_master.address
		.fpga_only_master_master_waitrequest                              (fpga_only_master_master_waitrequest),                              //                                                           .waitrequest
		.fpga_only_master_master_byteenable                               (fpga_only_master_master_byteenable),                               //                                                           .byteenable
		.fpga_only_master_master_read                                     (fpga_only_master_master_read),                                     //                                                           .read
		.fpga_only_master_master_readdata                                 (fpga_only_master_master_readdata),                                 //                                                           .readdata
		.fpga_only_master_master_readdatavalid                            (fpga_only_master_master_readdatavalid),                            //                                                           .readdatavalid
		.fpga_only_master_master_write                                    (fpga_only_master_master_write),                                    //                                                           .write
		.fpga_only_master_master_writedata                                (fpga_only_master_master_writedata),                                //                                                           .writedata
		.I2C_avalon_bridge_0_avalon_slave_0_address                       (mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_address),     //                         I2C_avalon_bridge_0_avalon_slave_0.address
		.I2C_avalon_bridge_0_avalon_slave_0_write                         (mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_write),       //                                                           .write
		.I2C_avalon_bridge_0_avalon_slave_0_read                          (mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_read),        //                                                           .read
		.I2C_avalon_bridge_0_avalon_slave_0_readdata                      (mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_readdata),    //                                                           .readdata
		.I2C_avalon_bridge_0_avalon_slave_0_writedata                     (mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_writedata),   //                                                           .writedata
		.I2C_avalon_bridge_0_avalon_slave_0_waitrequest                   (mm_interconnect_0_i2c_avalon_bridge_0_avalon_slave_0_waitrequest), //                                                           .waitrequest
		.I2C_avalon_bridge_1_avalon_slave_0_address                       (mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_address),     //                         I2C_avalon_bridge_1_avalon_slave_0.address
		.I2C_avalon_bridge_1_avalon_slave_0_write                         (mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_write),       //                                                           .write
		.I2C_avalon_bridge_1_avalon_slave_0_read                          (mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_read),        //                                                           .read
		.I2C_avalon_bridge_1_avalon_slave_0_readdata                      (mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_readdata),    //                                                           .readdata
		.I2C_avalon_bridge_1_avalon_slave_0_writedata                     (mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_writedata),   //                                                           .writedata
		.I2C_avalon_bridge_1_avalon_slave_0_waitrequest                   (mm_interconnect_0_i2c_avalon_bridge_1_avalon_slave_0_waitrequest), //                                                           .waitrequest
		.intr_capturer_0_avalon_slave_0_address                           (mm_interconnect_0_intr_capturer_0_avalon_slave_0_address),         //                             intr_capturer_0_avalon_slave_0.address
		.intr_capturer_0_avalon_slave_0_read                              (mm_interconnect_0_intr_capturer_0_avalon_slave_0_read),            //                                                           .read
		.intr_capturer_0_avalon_slave_0_readdata                          (mm_interconnect_0_intr_capturer_0_avalon_slave_0_readdata),        //                                                           .readdata
		.jtag_uart_avalon_jtag_slave_address                              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),            //                                jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),              //                                                           .write
		.jtag_uart_avalon_jtag_slave_read                                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),               //                                                           .read
		.jtag_uart_avalon_jtag_slave_readdata                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),           //                                                           .readdata
		.jtag_uart_avalon_jtag_slave_writedata                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),          //                                                           .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),        //                                                           .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),         //                                                           .chipselect
		.onchip_memory2_0_s1_address                                      (mm_interconnect_0_onchip_memory2_0_s1_address),                    //                                        onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                        (mm_interconnect_0_onchip_memory2_0_s1_write),                      //                                                           .write
		.onchip_memory2_0_s1_readdata                                     (mm_interconnect_0_onchip_memory2_0_s1_readdata),                   //                                                           .readdata
		.onchip_memory2_0_s1_writedata                                    (mm_interconnect_0_onchip_memory2_0_s1_writedata),                  //                                                           .writedata
		.onchip_memory2_0_s1_byteenable                                   (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                 //                                                           .byteenable
		.onchip_memory2_0_s1_chipselect                                   (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                 //                                                           .chipselect
		.onchip_memory2_0_s1_clken                                        (mm_interconnect_0_onchip_memory2_0_s1_clken),                      //                                                           .clken
		.sysid_qsys_control_slave_address                                 (mm_interconnect_0_sysid_qsys_control_slave_address),               //                                   sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                                (mm_interconnect_0_sysid_qsys_control_slave_readdata)               //                                                           .readdata
	);

	soc_system_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_f2h_axi_slave_awid                                            (mm_interconnect_1_hps_0_f2h_axi_slave_awid),    //                                           hps_0_f2h_axi_slave.awid
		.hps_0_f2h_axi_slave_awaddr                                          (mm_interconnect_1_hps_0_f2h_axi_slave_awaddr),  //                                                              .awaddr
		.hps_0_f2h_axi_slave_awlen                                           (mm_interconnect_1_hps_0_f2h_axi_slave_awlen),   //                                                              .awlen
		.hps_0_f2h_axi_slave_awsize                                          (mm_interconnect_1_hps_0_f2h_axi_slave_awsize),  //                                                              .awsize
		.hps_0_f2h_axi_slave_awburst                                         (mm_interconnect_1_hps_0_f2h_axi_slave_awburst), //                                                              .awburst
		.hps_0_f2h_axi_slave_awlock                                          (mm_interconnect_1_hps_0_f2h_axi_slave_awlock),  //                                                              .awlock
		.hps_0_f2h_axi_slave_awcache                                         (mm_interconnect_1_hps_0_f2h_axi_slave_awcache), //                                                              .awcache
		.hps_0_f2h_axi_slave_awprot                                          (mm_interconnect_1_hps_0_f2h_axi_slave_awprot),  //                                                              .awprot
		.hps_0_f2h_axi_slave_awuser                                          (mm_interconnect_1_hps_0_f2h_axi_slave_awuser),  //                                                              .awuser
		.hps_0_f2h_axi_slave_awvalid                                         (mm_interconnect_1_hps_0_f2h_axi_slave_awvalid), //                                                              .awvalid
		.hps_0_f2h_axi_slave_awready                                         (mm_interconnect_1_hps_0_f2h_axi_slave_awready), //                                                              .awready
		.hps_0_f2h_axi_slave_wid                                             (mm_interconnect_1_hps_0_f2h_axi_slave_wid),     //                                                              .wid
		.hps_0_f2h_axi_slave_wdata                                           (mm_interconnect_1_hps_0_f2h_axi_slave_wdata),   //                                                              .wdata
		.hps_0_f2h_axi_slave_wstrb                                           (mm_interconnect_1_hps_0_f2h_axi_slave_wstrb),   //                                                              .wstrb
		.hps_0_f2h_axi_slave_wlast                                           (mm_interconnect_1_hps_0_f2h_axi_slave_wlast),   //                                                              .wlast
		.hps_0_f2h_axi_slave_wvalid                                          (mm_interconnect_1_hps_0_f2h_axi_slave_wvalid),  //                                                              .wvalid
		.hps_0_f2h_axi_slave_wready                                          (mm_interconnect_1_hps_0_f2h_axi_slave_wready),  //                                                              .wready
		.hps_0_f2h_axi_slave_bid                                             (mm_interconnect_1_hps_0_f2h_axi_slave_bid),     //                                                              .bid
		.hps_0_f2h_axi_slave_bresp                                           (mm_interconnect_1_hps_0_f2h_axi_slave_bresp),   //                                                              .bresp
		.hps_0_f2h_axi_slave_bvalid                                          (mm_interconnect_1_hps_0_f2h_axi_slave_bvalid),  //                                                              .bvalid
		.hps_0_f2h_axi_slave_bready                                          (mm_interconnect_1_hps_0_f2h_axi_slave_bready),  //                                                              .bready
		.hps_0_f2h_axi_slave_arid                                            (mm_interconnect_1_hps_0_f2h_axi_slave_arid),    //                                                              .arid
		.hps_0_f2h_axi_slave_araddr                                          (mm_interconnect_1_hps_0_f2h_axi_slave_araddr),  //                                                              .araddr
		.hps_0_f2h_axi_slave_arlen                                           (mm_interconnect_1_hps_0_f2h_axi_slave_arlen),   //                                                              .arlen
		.hps_0_f2h_axi_slave_arsize                                          (mm_interconnect_1_hps_0_f2h_axi_slave_arsize),  //                                                              .arsize
		.hps_0_f2h_axi_slave_arburst                                         (mm_interconnect_1_hps_0_f2h_axi_slave_arburst), //                                                              .arburst
		.hps_0_f2h_axi_slave_arlock                                          (mm_interconnect_1_hps_0_f2h_axi_slave_arlock),  //                                                              .arlock
		.hps_0_f2h_axi_slave_arcache                                         (mm_interconnect_1_hps_0_f2h_axi_slave_arcache), //                                                              .arcache
		.hps_0_f2h_axi_slave_arprot                                          (mm_interconnect_1_hps_0_f2h_axi_slave_arprot),  //                                                              .arprot
		.hps_0_f2h_axi_slave_aruser                                          (mm_interconnect_1_hps_0_f2h_axi_slave_aruser),  //                                                              .aruser
		.hps_0_f2h_axi_slave_arvalid                                         (mm_interconnect_1_hps_0_f2h_axi_slave_arvalid), //                                                              .arvalid
		.hps_0_f2h_axi_slave_arready                                         (mm_interconnect_1_hps_0_f2h_axi_slave_arready), //                                                              .arready
		.hps_0_f2h_axi_slave_rid                                             (mm_interconnect_1_hps_0_f2h_axi_slave_rid),     //                                                              .rid
		.hps_0_f2h_axi_slave_rdata                                           (mm_interconnect_1_hps_0_f2h_axi_slave_rdata),   //                                                              .rdata
		.hps_0_f2h_axi_slave_rresp                                           (mm_interconnect_1_hps_0_f2h_axi_slave_rresp),   //                                                              .rresp
		.hps_0_f2h_axi_slave_rlast                                           (mm_interconnect_1_hps_0_f2h_axi_slave_rlast),   //                                                              .rlast
		.hps_0_f2h_axi_slave_rvalid                                          (mm_interconnect_1_hps_0_f2h_axi_slave_rvalid),  //                                                              .rvalid
		.hps_0_f2h_axi_slave_rready                                          (mm_interconnect_1_hps_0_f2h_axi_slave_rready),  //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                       //                                                     clk_0_clk.clk
		.hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset    (rst_controller_001_reset_out_reset),            //    hps_0_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
		.hps_only_master_clk_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                //               hps_only_master_clk_reset_reset_bridge_in_reset.reset
		.hps_only_master_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                // hps_only_master_master_translator_reset_reset_bridge_in_reset.reset
		.hps_only_master_master_address                                      (hps_only_master_master_address),                //                                        hps_only_master_master.address
		.hps_only_master_master_waitrequest                                  (hps_only_master_master_waitrequest),            //                                                              .waitrequest
		.hps_only_master_master_byteenable                                   (hps_only_master_master_byteenable),             //                                                              .byteenable
		.hps_only_master_master_read                                         (hps_only_master_master_read),                   //                                                              .read
		.hps_only_master_master_readdata                                     (hps_only_master_master_readdata),               //                                                              .readdata
		.hps_only_master_master_readdatavalid                                (hps_only_master_master_readdatavalid),          //                                                              .readdatavalid
		.hps_only_master_master_write                                        (hps_only_master_master_write),                  //                                                              .write
		.hps_only_master_master_writedata                                    (hps_only_master_master_writedata)               //                                                              .writedata
	);

	soc_system_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	soc_system_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_002 (
		.clk           (clk_clk),                                //       clk.clk
		.reset         (rst_controller_reset_out_reset),         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),               // receiver0.irq
		.sender_irq    (intr_capturer_0_interrupt_receiver_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
